module docker

import io

struct ChunkedResponseStream {
	reader io.Reader
}


