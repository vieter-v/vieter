module cron

import cli
import vieter_v.conf as vconf

struct Config {
pub:
	log_level               string = 'WARN'
	api_key                 string
	address                 string
	data_dir                string
	base_image              string = 'archlinux:base-devel'
	max_concurrent_builds   int    = 1
	api_update_frequency    int    = 15
	image_rebuild_frequency int    = 1440
	// Replicates the behavior of the original cron system
	global_schedule string = '0 3'
}

// cmd returns the cli module that handles the cron daemon.
pub fn cmd() cli.Command {
	return cli.Command{
		name: 'cron'
		description: 'Start the cron service that periodically runs builds.'
		execute: fn (cmd cli.Command) ? {
			config_file := cmd.flags.get_string('config-file')?
			conf := vconf.load<Config>(prefix: 'VIETER_', default_path: config_file)?

			cron(conf)?
		}
	}
}
