module git

pub struct GitRepo {
pub:
	url    string [required]
	branch string [required]
}
