module console
